library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity top is
    port (
        clk   : in std_logic
    );
end entity;

architecture behavourial of top is

begin

end architecture;