library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library vunit_lib;
context vunit_lib.vunit_context;

entity tb_top is
  generic (runner_cfg : string);
end entity;

architecture tb of tb_top is
begin

end architecture;